data:http://ns.logic.ly/1.6;base64,tVtdcxy5kfwrCjrCT4MWqlCFKvgsx/m8L36w/XBxD/d00R9oLy+4pGJ3FNb+eyemR7ujIbvdY1KxCkoaDTmJQlZmFtD7+4env9+PDz+/+/zDw+NPH+6+Px4//u79+8efutM/dA8/v6cu3/3h90/D/9fx+O7488f64e6hH+rDf355x927T/fTh7uc+mmswxQiOQeRKGFwlkCxkuZSMtf+7t3nD3eBuCtmJYlpjFFTuXv384c7Zes0ZSfORl6I7979+HTsj/dPjx/u4t27Y/18/HD3p++f7sd69/4K0U//uD+O319D4sTsRfvQ4+cC0tiH0nsfbPQ6xFhLidMJksSOc2EVvN1TUlkQkXVFtRSOhTyWa0RPn44fPx1Rtbl/+Ok5pqcfr/EMJZH1lAPPNQZJQwplSilUolqtVKl5OOEpRJ0lV805eyZbKkROHRAmKiwZf/ErPPePCxx5BqV/nK6xyKheR6KQxClI5CGUcbIwTBMqkSKn9qnAQtGsy9i+XEyMqegZTMIuckR9I8fEbitoeOdmGYqSQJXg0eYgmS14kRqGQammVI00ngAljl12MEQ1GnDm826VzpXxbZycE4nLbdv1MqqYxSdFXSgzUI0yhYGGARQqIEROYLZtoSLAKpE1m7ooivYWoDT5OPXuIUtRgOIaPM0UfB7Zsw+jG22B4gZKGa+VFD0qvQWoibjMlUuweTCAKlPoB5pDmkca1SQVGhdQVDpCRZK2Nsd3nTAl5Y48RwHjDQu8sVAvMLxaRc1LH4TmHGQ2DkXrFHygiWlMI5At3Q8qo5Im4BuRkNgJUaN9xt6Zu1BM10X6wu+0B8s4RQJl0PnjgB3jQUKB/oToA5p5Fu+ZT1iyaCfqxRJ2xpkWKAws4HZ0MohUpnjN7ZvA9FLmNIE0OoxTkL7mgI4HfSaP/VzHeRwXpVaVDqs3NBMEvDQBbJQ27SDP0KWYIdZJ1jp/F5hhyGJT8QDiAkwEjQepQ8iVKoo/Ow9Lg5mULqOdskDU3WJaaGMJSon9EXhHTrwfy8ss9im6FR9CHKVgo2LToyEHkuqsPEzYhEUWs4PF0JqSYS5wrKW1RLhzNkrgcFZw6U1UiGiy2FMKI7wRfGZGrw+Ev8aYSqm9ZdtCpeAPw8miSjm33C2gHp+OzxDNtY+qHvrmZ5Jgsh4z6mR57tXGcegXQsNNu5wKPpggldF4YbRG2EcWdIU1WiuvMZr2oJl0JhhpDNPI6Pcxz6GIwNsozzNkpu/lrD0mXQEkCE/KRMVPYIADGFEzhUQbemE3lof7v39//L/h08PwTKNnm1CQGYaKTARaABLP8NfRezBMYeKLnRHj04ujhILWdkt56TKGKMFiIkQgNf/4GtMzIC9FshJh8VM/BVg9zKtQQW/1pYWzHp5dkve6YEjorcKAhWThyGoLl9U6Sg6+5LZT6vnFSPbf8be/+fzH/9gHqdfsNU41iA6IZFhcGOZ5DlGqNIkZhvncX4KwE1EFMMrIXBbxUXc4mhlLU0JP10w+Q3php15Cw3ka01CGMFbsFFQOmWOUPkzAVeHazUlPaLh4hyaCh0FjnH0pkDG0pyABZQB1eSaEC5g/3lCemOaSZxlDKrAIaBpMVKuFPE6FpjmPOaUzoNJ0hiPsXUEaP0tz6uAaCjeLSZ5pz4Lnv/ZBGVkmGnoK5qk2AjN2SucAeHWwOdk0TxtQEBc7ReygplBRkd5ezvM3FAdhywYpY4C8gsQpItgjWARLoId5L9zLBiLoccdsouhxyYhDL5fnu73JcJprTWPGvNOjPn0fUZ9hxJfUI8HWpGP6Je+AHwUaCK2jtORni9IR5K/FC43w1ysw9fPHpx+Pf+1/AIDv+mP/L0V6ZSgjygoTiwPUUeYI4xjMwgS1Gysom+si02y5S9kMBgIhiEILSMooJDIZdBMivkKoE7wdVg8KyzxICv0c0W0V4w+GLQpzGqesPcogS2xFMG0JQzkyRgzY+0LuyNSlNpAheDA97/2b5p889HMPlwxaoUEyYw+ROxERMRghH0J0daE3yNYhvIJumLzaXHQC48wd9hPhByKP5ljLHbuwOOVhwoLCJCOoZFMOXltSHSMCPT5BdLEv5K0OOwWlNpRH86KJGFwxOWN0tZyjaV6z0l1YxgpF9CEivOOLkGJGdQXL5ziOEyRoKItAw7Q7tB3CYQJBSi5nSQSPirV5QyD18brr17GsW6lPLCnzFDIaC6I4RYRF5MRaBXDGISuPX0bV3KECiBmKkQfz82LvRhgNCxTBqUAq8r+w0lUgbUpGCkNZBmme3ivmd+JAaD2eINlWroAgOTdnt2WjDOlMJBkCJnotiv+7QFIsA2JWH6wfMU70Y4ESwjBmEGaSeWwT8BYQb86l0no6IXvpvw2kopV50gHZZkoAwh7KaBowv2Fkbw7iv1TEuxhhl8IEIclLDETk6toxELQa+YKuD312RD+zWSHFFLDfCBSzV2DpGZUBOTgiUeQFAcSkAyPxaY65IpOfLRP8RYWssQYSrWmNsTsjRR0xW1I7JsBggyjahqs6MyKF29C37uS6VASRAWZNEW1cSizn3AeEbTpuIxess/j1Ic8iuf+7NwEKTzMyVTADWTEMQ3wd22VDneGAc9QynFOoa9fUzBnBGYFzkbkWDBF61BCWpTDzyxHwb5+OO6uT0jgm6yGzyFrihHwDIcFgPqAQUx55jF+qg0iKOA7PQFgGuoW4GNWhutjBCMlJfD2Un6vz/MzpRTSSsUlIBCBuBHeGIkAzDVC9kmrNqU72Za8SIf8heMIEYEN2zn9WuhYIUUXDWmgFzU7mEH74NI8eMJqgNpMWOBKMcmoHPNTn6XQCuY4GGDrO7GA2fiGlvozm+ST8clCv2oZdzFAjcpbYjLCFlxBMM5JWckVOXsy6BT1HFyGkc2PJCUxgDDWY1iUKt2OMUwh7Ac5fPj0c7z8+1M/1x324vE6TZdZgXBAiiNDvGDeD6cCz5gojPJ+ktH5Hs8MTKZucj5monV6A3ykik1qE8rwcaeoPXwMbnx4fgQzvOuew//nzd3sPmJdv+PPjVD//qiin7993CHt6/6/f/vHp/rEJUogd/h2ZsmQMjdqcTQ/hdIweE+QUPYL0zYdyYikGKMea8Zosb4LqtwMm8uKR15e471h2fYn7TuG+XuIqmH2nsetg9p187QSz7xR2Hcy+M8GdYPadvq6D2XcMtxPMvnuOt2wL2gCza2Ubldm1mEsw6dce9dzMPCLbW4beeDpslG0fId4SKV8gZdhtm6oI9YZ28CEevn7N/RCcutiOaRKXVJr0ra9mX6+95Wo2SLBPhd4SzIVQYxSBQ1pBqkgY05KhtKfrjtjUWBMEOMkWMfYdSq+j33dYu4I+HpTgmBjnpBhyeoSTryLdd1C9jnTfQe6GIXI7QcXkCcVLcHg+aOpIWrpvNyqpDerr4HeV6S2tji7LjI1Fd0m7KUet2VCxDb3fVai3xMpXyaMUDAXtuBhYkS4QKqTd60ekEWT2iIH721X6dh//utKIbZ1BxkAKJGaxDeV4be/d7vIXUDlHMALJzTWhlwT2cbh+jQ4oG15CtJOEFN5O8b/dcm7PCZfLKdquGbwpIUoPZzycQ6xw2wX4Ssk5H9r7CpOoSjvLKXwI7WC7XRAI+rpNot9Qg24n10VroC86FUhPZDf8l9uOXb1mIGBBq7tJljZVY977dp1+OwH5615pN5oYuCICQOSsG73y2srfTq6NyusLlQffQL0OI39p19oY2oRkfT37cuj6evbdAe6dfXbdN2xY667T9y3FxzAdFQGgUBIqh9SGSHA4Srbsm0Pka7HvOyBf5TC6t0MiKIZWMwTZDQq/Fum+a4VVpO1MEAkG7l8yZlza8NDXIt130L+KNHGnEG4sNWqClOWNPtr3URvbv+sCYC19l9wJ9qDI6RAc6RBu0sX2gEZ0CCm0jTeou29DN2bZXXcGK9jbtXOG7SWj3B5NSvkQcuft1Ad/Pt1i6kZI3Nc269j3XTOsYE+nS1gS0WgE72gJsVPipMkRVdojMhuU2adWG/l218XECnSNuY25hhzSHkUriFjYBwQsasOaJ/zaYMyrDfvmxvwqYlGH6QFUz7B9/H5KWIiFDuDtiMzJkh7a27InhQkVF49FDyV2bbK31hntVm8jRL42vt++wovNkdOTQwgiGTtZpLVzW2HUcnqQCHoEjm3Fw1eCv13hL5si0mnwaBiTlOhbY/9r49TtSC+IBLnpSsztGrc9gWP6JatrJCqW2pFiET0AFgZswc8yIdDGEN8lNm9Qbbf3uaRvOF3dHgwu1VVbOkSnOFBm+O0prD9/UTIG2zaXx3K61f6GvX/7er4abBlN3HT19IgbR9lA+uqTmpvj5KVKWXtwqkB41PEV3GmVbxcXGAPR1xgC25HjARzrqD1DhPkQ4rWV1V/LpNvXc8mk5B0AtvvjdrNflqnv+jX8oXNiKQp4UICNoe+1F0v7bsVXT/wyadeAtlM0jD4bKXTfB71l2S9O10GKLsGWYVfOAm/bUtPXIr29NS+Qwqq69siOebsn5u17gNcivV33L5DCUBE5TdthdWYB5MVfNUdMyxkd6e35gG+H/vZwcIEetoPpXpsGRkyp8Vzn9+f/zekP/wQ=